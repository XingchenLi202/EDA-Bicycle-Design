module ecode(clock,a,b);
input [3:0] a;
input clock;
output [7:0] b;
reg [7:0] b;

always@(posedge clock)
	begin
	  
		case (a)
			4'b0000: b = 8'b00111111;//1000000; // 0
			4'b0001: b = 8'b00000110;//1111001; // 1
			4'b0010: b = 8'b01011011;//0100100; // 2
			4'b0011: b = 8'b01001111;//0110000; // 3
			4'b0100: b = 8'b01100110;//0011001; // 4
			4'b0101: b = 8'b01101101;//0010010; // 5
			4'b0110: b = 8'b01111101;//0000010; // 6
			4'b0111: b = 8'b00000111;//1111000; // 7
			4'b1000: b = 8'b01111111;//0000000; // 8
			4'b1001: b = 8'b01101111;//0010000; // 9
			default  b = 8'b00111111;//1000000; // 0
		endcase
	end
endmodule